library ieee;
use